library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.PIPECPU_STD.ALL;

entity pipeCPU is
  port(
        clk : in std_logic;
        rst : in std_logic;

        -- KEYBOARD --
        PS2KeyboardCLK : in std_logic;
        PS2KeyboardData : in std_logic;
        
        -- VGA ENGINE --
        vga_r  : out std_logic_vector(2 downto 0);
        vga_g  : out std_logic_vector(2 downto 0);
        vga_b  : out std_logic_vector(2 downto 1);
        h_sync : out std_logic;
        v_sync : out std_logic

  );
end pipeCPU;

architecture Behavioral of pipeCPU is
  -------------------------- CONSTANTS ----------------------------
  constant NOP : unsigned(31 downto 0) := (others => 0); -- NOP variabl
  
  ----------------------- INTERNAL SIGNALS ------------------------
  signal IR1 IR2, IR3, IR4 : unsigned(31 downto 0);
  signal IR1_next, IR2_next, IR3_next, IR4_next : unsigned(31 downto 0);
  signal pm_out : in unsigned(31 downto 0);
  signal pipe_control_signal : in unsigned(1 downto 0);

  -------------------------- ALIASES ------------------------------
  
  ---------------------- EXTERNAL COMPONENTS ------------------------
  --- VGA ENGINE ---
  component vga_engine is
  port (
        clk		 : in std_logic;
        rst    : in std_logic;
        
        char	   : in  unsigned(7 downto 0);
        fg_color : in  unsigned(7 downto 0);
        bg_color : in  unsigned(7 downto 0);
        addr	   : out unsigned(15 downto 0);
        
        vga_r  : out std_logic_vector(2 downto 0);
        vga_g  : out std_logic_vector(2 downto 0);
        vga_b  : out std_logic_vector(2 downto 1);
        h_sync : out std_logic;
        v_sync : out std_logic
       );
  end component;
  


  ---------------------- INTERNAL COMPONENTS ------------------------

  ----------- ControlUnit ------------
  component control_unit is
  port (
        clk : in std_logic;
        rst : in std_logic;
        -- IR in
        IR1 : in unsigned(31 downto 0);
        IR2 : in unsigned(31 downto 0);
        IR3 : in unsigned(31 downto 0);
        IR4 : in unsigned(31 downto 0);
        -- Flags input
        Z_flag : in std_logic;
        N_flag : in std_logic;
        O_flag : in std_logic;
        C_flag : in std_logic;
        -- Pipeline
        pipe_control_signal : out unsigned(1 downto 0);        
        -- PM 
        pm_control_signal : out unsigned(2 downto 0);
        -- RegisterFile control SIGNALS
        rf_read_d_or_b_control_signal : out std_logic;
        rf_write_d_control_signal : out std_logic;
        -- DataForwarding        
        df_control_signal : out unsigned(5 downto 0);
        -- ALU control signals  
        alu_update_flags_control_signal : out std_logic; -- 1 for true 0 for false
        alu_data_size_control_signal : out byte_mode;
        alu_op_control_signal : out op_code;
        -- KEYBOARD
        keyboard_read_signal : out std_logic;        
        -- DataMemory
        dm_write_or_read_control_signal : out std_logic;
        dm_size_mode_control_signal : out byte_mode;
        -- VideoMemory
        vm_write_enable_control_signal : out std_logic;
        -- WriteBackLogic
        wb_control_signal : out unsigned(1 downto 0)
  );


  ----------- ALU ------------
  component ALU is
  port (
        clk : in std_logic;
        rst : in std_logic;
        
        update_flags_control_signal : in unsigned(0 downto 0);
        data_size_control_signal : in byte_mode;
        alu_op_control_signal : in unsigned(5 downto 0);

        alu_a : in unsigned(31 downto 0); -- rA
        alu_b : in unsigned(31 downto 0); -- rB or IMM

        alu_res : out unsigned(31 downto 0);

        Z_flag, N_flag, O_flag, C_flag : buffer std_logic
  );
  
  ------- VIDEO MEMORY -------
  component video_memory is
  port (
        clk : in std_logic;
        rst : in std_logic;
        
        -- User port
        write_address : in unsigned(15 downto 0);
        write_data    : in unsigned(15 downto 0);
        write_enable  : in std_logic; -- Should write if true

        -- VGA engine port
        read_address : in  unsigned(15 downto 0);
        char         : out unsigned(7 downto 0);
        fg_color     : out unsigned(7 downto 0);
        bg_color     : out unsigned(7 downto 0)
       );
  end component;  


  ------------------------ MAPPING SIGNALS -----------------------
  signal map_update_flags_control_signal : std_logic;
  signal map_data_size_control_signal : byte_mode;
  signal map_alu_op_control_signal : unsigned(5 downto 0);
  signal map_alu_a : unsigned(31 downto 0);
  signal map_alu_b : unsigned(31 downto 0);
  signal map_alu_res : unsigned(31 downto 0);
  signal map_Z_flag, map_N_flag, map_O_flag, map_C_flag : buffer std_logic;
  
  signal map_vm_write_addres : unsigned(15 downto 0);
  signal map_vm_write_data : unsigned(15 downto 0);
  signal map_vm_write_enable_control_signal : std_logic;
  
  signal map_vga_address : unsigned(15 downto 0);
  signal map_vga_char : unsigned(7 downto 0);
  signal map_vga_fg_color : unsigned(7 downto 0);
  signal map_vga_bg_color : unsigned(7 downto 0);

begin

  ------------------------- PORT MAPPINGS ------------------------
  
  ----------- ControlUnit ------------
 -- u_control_unit : control_unit
  --port map (
    --alu_update_flags_control_signal => map_update_flags_control_signal, -- OUT

  ----------- ALU ------------
  U_ALU : ALU
  port map (
    clk => clk,                                                     -- IN
    rst => rst,                                                     -- IN
    update_flags_control_signal => map_update_flags_control_signal, -- IN
    data_size_control_signal => map_data_size_control_signal,       -- IN
    alu_op_control_signal => map_alu_op_control_signal,             -- IN
    alu_a => map_alu_a,                                             -- IN
    alu_b => map_alu_b,                                             -- IN

    alu_res => map_alu_res,                                         -- OUT
    Z_flag => map_Z_flag,                                           -- OUT
    N_flag => map_N_flag,                                           -- OUT
    O_flag => map_O_flag,                                           -- OUT
    C_flag => map_C_flag                                            -- OUT
  );


   U_VGA : vga_engine port map (
    -- INTERNAL
    clk => clk,                        -- IN
    rst => rst,                        -- IN
    char => map_vga_char,              -- IN
    fg_color => map_vga_fg_color,      -- IN
    bg_color => map_vga_bg_color,      -- IN
    addr => map_vga_address,           -- OUT
    -- EXTERNAL
    vga_r => vga_r,                    -- OUT
    vga_g => vga_g,                    -- OUT
    vga_b => vga_b,                    -- OUT
    h_sync => h_sync,                  -- OUT
    v_sync => v_sync                   -- OUT
   );



  -------------------------- INTERNAL LOGIC ----------------------------

  -- Data stall / jump mux logic
  with pipe_control_signals select
  IR1_next <= NOP when PIPE_JMP,
              IR1 when PIPE_STALL,
              pm_out when others;
    
  with pipe_control_signals select
  IR2_next <= NOP when PIPE_STALL,
              IR1 when others;
  
  IR3_next <= IR2;

  IR4_next <= IR3;

  -- Update registers on clock cycle
  process(clk)
  begin
    if rising_edge(clk) then 
      if rst = '1' then 
        IR1 <= NOP;
        IR2 <= NOP;
        IR3 <= NOP;
        IR4 <= NOP;
      else
        IR1 <= IR1_next;
        IR2 <= IR2_next;
        IR3 <= IR3_next;
        IR4 <= IR4_next;
      end if;
    end if;
  

  --------------------------------- END -------------------------------
  end;

end architecture;    

