library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.PIPECPU_STD.ALL;

package data_file is
  
  constant data0 : data_chunk_array := (
--$DATA1
X"20",
X"20",
X"20",
X"2d",
X"20",
X"20",
X"26",
X"20",
X"2d",
X"20",
X"20",
X"2f",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"26",
X"26",
X"20",
X"40",
X"40",
X"20",
X"40",
X"20",
X"26",
X"0a",
X"7c",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"40",
X"2a",
X"20",
X"20",
X"20",
X"40",
X"40",
X"40",
X"40",
X"20",
X"5e",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"40",
X"20",
X"20",
X"20",
X"26",
X"20",
X"40",
X"40",
X"20",
X"40",
X"20",
X"40",
X"0a",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"2f",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"40",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"00",
X"00",
X"92",
X"e0",
X"fc",
X"1c",
X"1f",
X"03",
X"e3",
X"fd",
X"2d",
X"4d",
X"24",
X"b6",
X"e9",
X"cf",
X"86",
X"06",
X"28",
X"00",
X"10",
X"80",
X"00",
X"00",
X"00",
X"73",
X"6c",
X"61",
X"78",
X"6e",
X"61",
X"6f",
X"63",
X"6e",
X"65",
X"6e",
X"5f",
X"6e",
X"00",
X"28",
X"05",
X"00",
X"00",
X"03",
X"02",
X"06",
X"53",
X"54",
X"2e",
X"00",
X"59",
X"58",
X"4e",
X"52",
X"20",
X"45",
X"4f",
X"41",
X"47",
X"0a",
X"4f",
X"41",
X"41",
X"52",
X"4b",
X"2e",
X"00",
X"44",
X"0a",
--$DATA1_END
others => X"00"
);
  constant data1 : data_chunk_array := (
--$DATA2
X"20",
X"20",
X"0a",
X"24",
X"20",
X"55",
X"2d",
X"0a",
X"24",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"3e",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"40",
X"40",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"25",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"7c",
X"7c",
X"20",
X"40",
X"40",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"40",
X"27",
X"2a",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"40",
X"20",
X"40",
X"26",
X"20",
X"40",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"27",
X"20",
X"20",
X"40",
X"40",
X"20",
X"40",
X"20",
X"2f",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"20",
X"40",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0f",
X"00",
X"00",
X"00",
X"02",
X"00",
X"00",
X"00",
X"63",
X"73",
X"74",
X"00",
X"67",
X"69",
X"77",
X"72",
X"73",
X"72",
X"61",
X"70",
X"74",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"03",
X"07",
X"54",
X"49",
X"2e",
X"50",
X"45",
X"20",
X"0a",
X"45",
X"45",
X"52",
X"20",
X"59",
X"41",
X"00",
X"4f",
X"41",
X"4c",
X"45",
X"49",
X"2e",
X"47",
X"42",
X"00",
--$DATA2_END
others => X"00"
);

  constant data2 : data_chunk_array := (
--$DATA3
X"20",
X"20",
X"20",
X"26",
X"20",
X"2d",
X"4f",
X"20",
X"26",
X"20",
X"20",
X"20",
X"00",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"40",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"2f",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"23",
X"26",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"40",
X"20",
X"20",
X"40",
X"26",
X"40",
X"40",
X"40",
X"20",
X"20",
X"20",
X"7e",
X"0a",
X"26",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"2e",
X"40",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"2a",
X"40",
X"26",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"40",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"26",
X"26",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"00",
X"49",
X"ff",
X"f0",
X"9c",
X"1e",
X"13",
X"83",
X"5f",
X"be",
X"6c",
X"cf",
X"76",
X"57",
X"41",
X"a6",
X"ea",
X"00",
X"1e",
X"00",
X"00",
X"e0",
X"00",
X"00",
X"64",
X"6f",
X"00",
X"72",
X"70",
X"00",
X"6e",
X"00",
X"65",
X"61",
X"00",
X"6b",
X"61",
X"00",
X"07",
X"1e",
X"01",
X"26",
X"02",
X"00",
X"04",
X"08",
X"41",
X"4e",
X"2e",
X"4c",
X"52",
X"57",
X"00",
X"53",
X"4e",
X"20",
X"50",
X"20",
X"49",
X"47",
X"4f",
X"41",
X"0a",
X"4d",
X"4e",
X"2e",
X"4f",
X"59",
--$DATA3_END
others => X"00"
);

  constant data3 : data_chunk_array := (
--$DATA4
X"24",
X"20",
X"4d",
X"20",
X"0a",
X"24",
X"53",
X"58",
X"20",
X"0a",
X"24",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"3e",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"40",
X"40",
X"20",
X"40",
X"3e",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"26",
X"20",
X"26",
X"20",
X"40",
X"26",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"7c",
X"40",
X"40",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"40",
X"2f",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"40",
X"20",
X"40",
X"20",
X"20",
X"20",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"20",
X"40",
X"40",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"20",
X"26",
X"20",
X"40",
X"3e",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"40",
X"3e",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"3e",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"20",
X"0a",
X"10",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"00",
X"00",
X"69",
X"00",
X"6d",
X"69",
X"6f",
X"72",
X"62",
X"73",
X"65",
X"76",
X"73",
X"65",
X"69",
X"0a",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"05",
X"00",
X"52",
X"47",
X"0a",
X"41",
X"20",
X"4f",
X"50",
X"53",
X"54",
X"54",
X"4c",
X"41",
X"4e",
X"4f",
X"4f",
X"41",
X"00",
X"41",
X"47",
X"0a",
X"4f",
X"45",
--$DATA4_END
others => X"00"
);
  
end data_file;
