library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library work;
use work.PIPECPU_STD.ALL;

entity control_unit is 

end control_unit;

architecture Behavioural of control_unit is 



end Behavioural;
