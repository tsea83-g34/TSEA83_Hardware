library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package CHARS is
  
  constant NUMBER_OF_CHARS : INTEGER := 128;
  constant CHAR_SIZE       : INTEGER := 16;
  constant CHAR_BIT_SIZE   : INTEGER := 4;
  
  type char_array is array (0 to NUMBER_OF_CHARS - 1) of UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0);
  
  -- ======== Chars ========
  
  constant CHARS : char_array := (

-- NULL_CHAR
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SOH
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- STX
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ETX
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EOT
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ENQ
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ACK
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- BEL
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- BS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- HT
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- LF
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- VT
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- FF
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- CR
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SO
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SI
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DLE
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DC1
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DC2
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DC3
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DC4
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- NAK
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SYN
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ETB
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- CAN
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EM
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SUB
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ESC
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- FS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- GS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- RS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- US
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SPACE
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EXCLAMATION_MARK
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DOUBLE_QUOTE
"0000000000000000" &
"0000011100111000" &
"0000011100111000" &
"0000011100111000" &
"0000011100111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- HASH
"0000000000000000" &
"0000000011000111" &
"0000000011000111" &
"0000000011000110" &
"0000000011000110" &
"0000111111111111" &
"0000000100001110" &
"0000000100001000" &
"0000000100001000" &
"0011111111111111" &
"0000011000111000" &
"0000011000110000" &
"0000111000110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DOLLAR
"0000000000000000" &
"0000000100000000" &
"0000111111110000" &
"0011100100110000" &
"0011100100000000" &
"1111100100000000" &
"0011111100000000" &
"0000111111110000" &
"0000000111111000" &
"0000000100111000" &
"0000000100111000" &
"0011000100111000" &
"0011111111110000" &
"0000000100000000" &
"0000000100000000" &
"0000000000000000",

-- PERCENT
"0000000000000000" &
"0000000000000000" &
"0000111100000000" &
"0011000011000000" &
"0011000011000000" &
"0011000011000000" &
"0000111100001110" &
"0000000111110000" &
"0000111000111110" &
"0000000011000001" &
"0000000011000001" &
"0000000011000001" &
"0000000000111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- AMPERSAND
"0000000000000000" &
"0000000111110000" &
"0000011000000000" &
"0000011000000000" &
"0000011000000000" &
"0000011100000000" &
"0000111100000000" &
"0000100011000111" &
"0011100011000111" &
"0011100000110111" &
"0011100000001110" &
"0000111000001110" &
"0000011111110111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SINGLE_QUOTE
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- LEFT_PARENTHESES
"0000000000000000" &
"0000000011110000" &
"0000000011000000" &
"0000000111000000" &
"0000000111000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000000111000000" &
"0000000111000000" &
"0000000011000000" &
"0000000011110000" &
"0000000000000000",

-- RIGHT_PARENTHESES
"0000000000000000" &
"0000011100000000" &
"0000000100000000" &
"0000000111000000" &
"0000000111000000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000111000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000000000000000",

-- STAR
"0000000000000000" &
"0000000100000000" &
"0011000100001000" &
"0000100100110000" &
"0000011111000000" &
"0000111111110000" &
"0011000100001000" &
"0000000100000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- PLUS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111111111110" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- COMMA
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000000000000000",

-- DASH
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- PERIOD
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SLASH
"0000000000000000" &
"0000000000001000" &
"0000000000111000" &
"0000000000110000" &
"0000000011110000" &
"0000000011000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000011000000000" &
"0000111000000000" &
"0000100000000000" &
"0011100000000000" &
"0011100000000000" &
"0000000000000000" &
"0000000000000000",

-- ZERO
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0000100000001000" &
"0011100000001110" &
"0011100000001110" &
"0011100111001110" &
"0011100111001110" &
"0011100000001110" &
"0011100000001110" &
"0000100000001000" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ONE
"0000000000000000" &
"0000111111000000" &
"0000111111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- TWO
"0000000000000000" &
"0011111111000000" &
"0011000011110000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000011110000" &
"0000000011110000" &
"0000000111000000" &
"0000011100000000" &
"0000111000000000" &
"0011100000000000" &
"0011111111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- THREE
"0000000000000000" &
"0000111111110000" &
"0000000000111110" &
"0000000000001110" &
"0000000000001110" &
"0000000000111000" &
"0000000111000000" &
"0000000000111000" &
"0000000000001110" &
"0000000000001110" &
"0000000000001110" &
"0011000000111000" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- FOUR
"0000000000000000" &
"0000000011111000" &
"0000000011111000" &
"0000000100111000" &
"0000000100111000" &
"0000011000111000" &
"0000111000111000" &
"0000100000111000" &
"0011100000111000" &
"0011111111111111" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- Five
"0000000000000000" &
"0000111111111000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111110000" &
"0000000000111000" &
"0000000000001110" &
"0000000000001110" &
"0000000000001110" &
"0000000000001110" &
"0011000000111000" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SIX
"0000000000000000" &
"0000011111111000" &
"0000111000000000" &
"0000111000000000" &
"0011100000000000" &
"0011100111110000" &
"0011111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SEVEN
"0000000000000000" &
"0011111111111000" &
"0000000000111000" &
"0000000000110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011000000" &
"0000000111000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EIGHT
"0000000000000000" &
"0000011111110000" &
"0011111000111110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- NINE
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111110" &
"0000011111001110" &
"0000000000001110" &
"0000000000111000" &
"0000000000111000" &
"0000111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- COLON
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SEMICOLON
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000000000000000",

-- LESS_THAN
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000111" &
"0000000000111110" &
"0000011111110000" &
"0011111000000000" &
"0011111000000000" &
"0000011111110000" &
"0000000000111111" &
"0000000000000110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EQUAL
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011111111111110" &
"0000000000000000" &
"0000000000000000" &
"0011111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- GREATER_THAN
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011000000000000" &
"0011111100000000" &
"0000000111110000" &
"0000000000001111" &
"0000000000111111" &
"0000000111110000" &
"0011111100000000" &
"0011000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- QUESTION_MARK
"0000000000000000" &
"0000111111110000" &
"0000100000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000011111000" &
"0000000111110000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- AT
"0000000000000000" &
"0000000000000000" &
"0000000111111000" &
"0000011000000110" &
"0000100000000001" &
"0011100011111111" &
"0011000111000111" &
"0011000100000001" &
"0011000100000001" &
"0011000111000111" &
"0011000011111111" &
"0000100000000000" &
"0000100000000000" &
"0000011100000000" &
"0000000111111110" &
"0000000000000000",

-- A
"0000000000000000" &
"0000000111000000" &
"0000011111000000" &
"0000011111110000" &
"0000011011110000" &
"0000011000110000" &
"0000111000110000" &
"0000111000111000" &
"0000100000111000" &
"0011111111111000" &
"0011100000001110" &
"0011000000001110" &
"1111000000000110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- B
"0000000000000000" &
"0011111111110000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011111111000000" &
"0011100000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000111110" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- C
"0000000000000000" &
"0000000111111110" &
"0000111000000110" &
"0000111000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0000111000000000" &
"0000111000000110" &
"0000000111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- D
"0000000000000000" &
"0011111111000000" &
"0011100000111000" &
"0011100000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000111000" &
"0011100000111000" &
"0011111111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- E
"0000000000000000" &
"0000111111111110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111111110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- F
"0000000000000000" &
"0000111111111110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111111110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- G
"0000000000000000" &
"0000000111111000" &
"0000111000001000" &
"0000111000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000111110" &
"0011100000001110" &
"0011100000001110" &
"0000100000001110" &
"0000111000001110" &
"0000000111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- H
"0000000000000000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011111111111110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- I
"0000000000000000" &
"0000111111111000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000111111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- J
"0000000000000000" &
"0000011111111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0011000011111000" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- K
"0000000000000000" &
"0011100000001110" &
"0011100000001000" &
"0011100000110000" &
"0011100011110000" &
"0011100111000000" &
"0011111111000000" &
"0011111011000000" &
"0011100011110000" &
"0011100000111000" &
"0011100000111000" &
"0011100000001110" &
"0011100000000111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- L
"0000000000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111111111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- M
"0000000000000000" &
"0011111000001111" &
"0011111000001111" &
"0011111000001111" &
"0011100100110111" &
"0011100100110111" &
"0011100100110111" &
"0011100011000111" &
"0011100011000111" &
"0011100000000111" &
"0011100000000111" &
"0011100000000111" &
"0011100000000111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- N
"0000000000000000" &
"0011111000001110" &
"0011111000001110" &
"0011111000001110" &
"0011111100001110" &
"0011100100001110" &
"0011100100001110" &
"0011100011001110" &
"0011100011001110" &
"0011100011111110" &
"0011100000111110" &
"0011100000111110" &
"0011100000111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- O
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- P
"0000000000000000" &
"0000111111111000" &
"0000111000001110" &
"0000111000000111" &
"0000111000000111" &
"0000111000000111" &
"0000111000001110" &
"0000111111111000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- Q
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001000" &
"0000111000111000" &
"0000011111110000" &
"0000000000111000" &
"0000000000001000" &
"0000000000000000",

-- R
"0000000000000000" &
"0011111111000000" &
"0011100011110000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100011110000" &
"0011111111000000" &
"0011100011110000" &
"0011100000110000" &
"0011100000001000" &
"0011100000001110" &
"0011100000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- S
"0000000000000000" &
"0000011111111000" &
"0000111000001000" &
"0011100000000000" &
"0011100000000000" &
"0011111000000000" &
"0000111111110000" &
"0000000111111000" &
"0000000000111110" &
"0000000000001110" &
"0000000000001110" &
"0011000000111000" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- T
"0000000000000000" &
"0011111111111111" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- U
"0000000000000000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- V
"0000000000000000" &
"0011000000001110" &
"0011000000001110" &
"0011100000001000" &
"0011100000001000" &
"0000100000111000" &
"0000100000111000" &
"0000111000110000" &
"0000011000110000" &
"0000011011110000" &
"0000011111110000" &
"0000011111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- W
"0000000000000000" &
"1111000000000111" &
"1111000000000110" &
"1111000000000110" &
"0011000111000110" &
"0011000111000110" &
"0011011111001110" &
"0011011011001110" &
"0011011011111110" &
"0011111000111000" &
"0011111000111000" &
"0000111000111000" &
"0000100000111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- X
"0000000000000000" &
"0011100000001110" &
"0000100000001000" &
"0000111000111000" &
"0000011000110000" &
"0000011111000000" &
"0000000111000000" &
"0000000111000000" &
"0000011111110000" &
"0000111000110000" &
"0000100000111000" &
"0011100000001110" &
"1111000000000110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- Y
"0000000000000000" &
"0011000000000110" &
"0011100000001110" &
"0000100000001000" &
"0000111000111000" &
"0000011111110000" &
"0000011111110000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- Z
"0000000000000000" &
"0011111111111110" &
"0000000000001110" &
"0000000000111000" &
"0000000000110000" &
"0000000011110000" &
"0000000111000000" &
"0000000111000000" &
"0000011100000000" &
"0000011000000000" &
"0000111000000000" &
"0011100000000000" &
"0011111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- LEFT_BRACKET
"0000000000000000" &
"0000000111111000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111111000" &
"0000000000000000",

-- BACK_SLASH
"0000000000000000" &
"0011100000000000" &
"0000100000000000" &
"0000100000000000" &
"0000111000000000" &
"0000011000000000" &
"0000011100000000" &
"0000000100000000" &
"0000000111000000" &
"0000000011000000" &
"0000000011110000" &
"0000000000110000" &
"0000000000111000" &
"0000000000001000" &
"0000000000000000" &
"0000000000000000",

-- RIGHT_BRACKET
"0000000000000000" &
"0000011111110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000011111110000" &
"0000000000000000",

-- HAT
"0000000000000000" &
"0000000111000000" &
"0000011111110000" &
"0000111000110000" &
"0011100000001000" &
"0011000000000110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- UNDERSCORE
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- LEFT_TICK
"0000011000000000" &
"0000011100000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- a_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111111110000" &
"0000100011111000" &
"0000000000111000" &
"0000000000111000" &
"0000111111111000" &
"0011100000111000" &
"0011100000111000" &
"0011100011111000" &
"0000111100111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- b_low
"0000000000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111011111000" &
"0000111100111000" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111100111000" &
"0000111011111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- c_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111111110" &
"0000011100000110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000011100000110" &
"0000000111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- d_low
"0000000000000000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000111100111000" &
"0000111011111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0000111011111000" &
"0000111100111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- e_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011111111111110" &
"0011100000000000" &
"0011100000000000" &
"0000111000000110" &
"0000011111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- f_low
"0000000000000000" &
"0000000011111110" &
"0000000111000000" &
"0000000111000000" &
"0000111111111110" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- g_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111100111000" &
"0000111011111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0000111011111000" &
"0000111100111000" &
"0000000000111000" &
"0000100011110000" &
"0000111111110000",

-- h_low
"0000000000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111011111000" &
"0000111100001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- i_low
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000111111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- j_low
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000111111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111100000000",

-- k_low
"0000000000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000001110" &
"0000111000111000" &
"0000111011110000" &
"0000111111000000" &
"0000111111110000" &
"0000111000111000" &
"0000111000001000" &
"0000111000001110" &
"0000111000000111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- l_low
"0000000000000000" &
"0000111111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000011111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- m_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011111100111000" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- n_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111011111000" &
"0000111100001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- o_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- p_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011100111110000" &
"0011111011110000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011111011110000" &
"0011100111110000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000",

-- q_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111100111000" &
"0000111011111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0000111011111000" &
"0000111100111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000",

-- r_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011100111110" &
"0000011111000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- s_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011111111000" &
"0000111000000000" &
"0000111000000000" &
"0000111100000000" &
"0000011111111000" &
"0000000000111110" &
"0000000000001110" &
"0000100000001110" &
"0000111111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- t_low
"0000000000000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0011111111111000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000000111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- u_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000111110" &
"0000011111001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- v_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011000000001110" &
"0011100000001000" &
"0000100000111000" &
"0000100000111000" &
"0000111000110000" &
"0000011011110000" &
"0000011011110000" &
"0000011111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- w_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"1111000000000111" &
"1111000000000110" &
"0011000000000110" &
"0011000111001110" &
"0011000111001110" &
"0011111011001000" &
"0011111011001000" &
"0000111000111000" &
"0000111000111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- x_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011100000001000" &
"0000111000111000" &
"0000011011110000" &
"0000011111000000" &
"0000000111000000" &
"0000011111000000" &
"0000111000110000" &
"0000100000111000" &
"0011100000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- y_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011000000001000" &
"0011000000111000" &
"0011100000111000" &
"0000100000110000" &
"0000111011110000" &
"0000011011000000" &
"0000011011000000" &
"0000011111000000" &
"0000000100000000" &
"0000011100000000" &
"0000011000000000" &
"0011111000000000",

-- z_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111111111110" &
"0000000000001110" &
"0000000000111000" &
"0000000011110000" &
"0000000011000000" &
"0000000111000000" &
"0000011100000000" &
"0000111000000000" &
"0000111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- CURLY_LEFT
"0000000000000000" &
"0000000011111000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000011111000",

-- PIPE
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000",

-- CURLY_RIGHT
"0000000000000000" &
"0011111100000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000111000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111100000000",

-- SWUNG_DASH
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111100000110" &
"0011000011111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DEL
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000"
);
  
  -- ======== Alias ========
  -- Indexes
  constant NULL_CHAR: INTEGER := 0;
  constant SOH: INTEGER := 1;
  constant STX: INTEGER := 2;
  constant ETX: INTEGER := 3;
  constant EOT: INTEGER := 4;
  constant ENQ: INTEGER := 5;
  constant ACK: INTEGER := 6;
  constant BEL: INTEGER := 7;
  constant BS: INTEGER := 8;
  constant HT: INTEGER := 9;
  constant LF: INTEGER := 10;
  constant VT: INTEGER := 11;
  constant FF: INTEGER := 12;
  constant CR: INTEGER := 13;
  constant SO: INTEGER := 14;
  constant SI: INTEGER := 15;
  constant DLE: INTEGER := 16;
  constant DC1: INTEGER := 17;
  constant DC2: INTEGER := 18;
  constant DC3: INTEGER := 19;
  constant DC4: INTEGER := 20;
  constant NAK: INTEGER := 21;
  constant SYN: INTEGER := 22;
  constant ETB: INTEGER := 23;
  constant CAN: INTEGER := 24;
  constant EM: INTEGER := 25;
  constant SUB: INTEGER := 26;
  constant ESC: INTEGER := 27;
  constant FS: INTEGER := 28;
  constant GS: INTEGER := 29;
  constant RS: INTEGER := 30;
  constant US: INTEGER := 31;
  constant SPACE: INTEGER := 32;
  constant EXCLAMATION_MARK: INTEGER := 33;
  constant DOUBLE_QUOTE: INTEGER := 34;
  constant HASH: INTEGER := 35;
  constant DOLLAR: INTEGER := 36;
  constant PERCENT: INTEGER := 37;
  constant AMPERSAND: INTEGER := 38;
  constant SINGLE_QUOTE: INTEGER := 39;
  constant LEFT_PARENTHESES: INTEGER := 40;
  constant RIGHT_PARENTHESES: INTEGER := 41;
  constant STAR: INTEGER := 42;
  constant PLUS: INTEGER := 43;
  constant COMMA: INTEGER := 44;
  constant DASH: INTEGER := 45;
  constant PERIOD: INTEGER := 46;
  constant SLASH: INTEGER := 47;
  constant ZERO: INTEGER := 48;
  constant ONE: INTEGER := 49;
  constant TWO: INTEGER := 50;
  constant THREE: INTEGER := 51;
  constant FOUR: INTEGER := 52;
  constant Five: INTEGER := 53;
  constant SIX: INTEGER := 54;
  constant SEVEN: INTEGER := 55;
  constant EIGHT: INTEGER := 56;
  constant NINE: INTEGER := 57;
  constant COLON: INTEGER := 58;
  constant SEMICOLON: INTEGER := 59;
  constant LESS_THAN: INTEGER := 60;
  constant EQUAL: INTEGER := 61;
  constant GREATER_THAN: INTEGER := 62;
  constant QUESTION_MARK: INTEGER := 63;
  constant AT: INTEGER := 64;
  constant A: INTEGER := 65;
  constant B: INTEGER := 66;
  constant C: INTEGER := 67;
  constant D: INTEGER := 68;
  constant E: INTEGER := 69;
  constant F: INTEGER := 70;
  constant G: INTEGER := 71;
  constant H: INTEGER := 72;
  constant I: INTEGER := 73;
  constant J: INTEGER := 74;
  constant K: INTEGER := 75;
  constant L: INTEGER := 76;
  constant M: INTEGER := 77;
  constant N: INTEGER := 78;
  constant O: INTEGER := 79;
  constant P: INTEGER := 80;
  constant Q: INTEGER := 81;
  constant R: INTEGER := 82;
  constant S: INTEGER := 83;
  constant T: INTEGER := 84;
  constant U: INTEGER := 85;
  constant V: INTEGER := 86;
  constant W: INTEGER := 87;
  constant X: INTEGER := 88;
  constant Y: INTEGER := 89;
  constant Z: INTEGER := 90;
  constant LEFT_BRACKET: INTEGER := 91;
  constant BACK_SLASH: INTEGER := 92;
  constant RIGHT_BRACKET: INTEGER := 93;
  constant HAT: INTEGER := 94;
  constant UNDERSCORE: INTEGER := 95;
  constant LEFT_TICK: INTEGER := 96;
  constant a_low: INTEGER := 97;
  constant b_low: INTEGER := 98;
  constant c_low: INTEGER := 99;
  constant d_low: INTEGER := 100;
  constant e_low: INTEGER := 101;
  constant f_low: INTEGER := 102;
  constant g_low: INTEGER := 103;
  constant h_low: INTEGER := 104;
  constant i_low: INTEGER := 105;
  constant j_low: INTEGER := 106;
  constant k_low: INTEGER := 107;
  constant l_low: INTEGER := 108;
  constant m_low: INTEGER := 109;
  constant n_low: INTEGER := 110;
  constant o_low: INTEGER := 111;
  constant p_low: INTEGER := 112;
  constant q_low: INTEGER := 113;
  constant r_low: INTEGER := 114;
  constant s_low: INTEGER := 115;
  constant t_low: INTEGER := 116;
  constant u_low: INTEGER := 117;
  constant v_low: INTEGER := 118;
  constant w_low: INTEGER := 119;
  constant x_low: INTEGER := 120;
  constant y_low: INTEGER := 121;
  constant z_low: INTEGER := 122;
  constant CURLY_LEFT: INTEGER := 123;
  constant PIPE: INTEGER := 124;
  constant CURLY_RIGHT: INTEGER := 125;
  constant SWUNG_DASH: INTEGER := 126;
  constant DEL: INTEGER := 127;

  -- Chars
  alias NULL_CHAR_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(0);
  alias SOH_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(1);
  alias STX_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(2);
  alias ETX_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(3);
  alias EOT_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(4);
  alias ENQ_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(5);
  alias ACK_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(6);
  alias BEL_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(7);
  alias BS_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(8);
  alias HT_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(9);
  alias LF_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(10);
  alias VT_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(11);
  alias FF_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(12);
  alias CR_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(13);
  alias SO_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(14);
  alias SI_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(15);
  alias DLE_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(16);
  alias DC1_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(17);
  alias DC2_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(18);
  alias DC3_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(19);
  alias DC4_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(20);
  alias NAK_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(21);
  alias SYN_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(22);
  alias ETB_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(23);
  alias CAN_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(24);
  alias EM_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(25);
  alias SUB_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(26);
  alias ESC_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(27);
  alias FS_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(28);
  alias GS_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(29);
  alias RS_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(30);
  alias US_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(31);
  alias SPACE_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(32);
  alias EXCLAMATION_MARK_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(33);
  alias DOUBLE_QUOTE_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(34);
  alias HASH_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(35);
  alias DOLLAR_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(36);
  alias PERCENT_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(37);
  alias AMPERSAND_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(38);
  alias SINGLE_QUOTE_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(39);
  alias LEFT_PARENTHESES_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(40);
  alias RIGHT_PARENTHESES_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(41);
  alias STAR_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(42);
  alias PLUS_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(43);
  alias COMMA_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(44);
  alias DASH_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(45);
  alias PERIOD_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(46);
  alias SLASH_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(47);
  alias ZERO_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(48);
  alias ONE_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(49);
  alias TWO_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(50);
  alias THREE_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(51);
  alias FOUR_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(52);
  alias Five_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(53);
  alias SIX_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(54);
  alias SEVEN_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(55);
  alias EIGHT_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(56);
  alias NINE_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(57);
  alias COLON_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(58);
  alias SEMICOLON_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(59);
  alias LESS_THAN_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(60);
  alias EQUAL_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(61);
  alias GREATER_THAN_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(62);
  alias QUESTION_MARK_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(63);
  alias AT_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(64);
  alias A_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(65);
  alias B_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(66);
  alias C_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(67);
  alias D_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(68);
  alias E_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(69);
  alias F_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(70);
  alias G_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(71);
  alias H_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(72);
  alias I_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(73);
  alias J_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(74);
  alias K_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(75);
  alias L_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(76);
  alias M_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(77);
  alias N_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(78);
  alias O_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(79);
  alias P_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(80);
  alias Q_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(81);
  alias R_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(82);
  alias S_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(83);
  alias T_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(84);
  alias U_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(85);
  alias V_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(86);
  alias W_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(87);
  alias X_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(88);
  alias Y_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(89);
  alias Z_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(90);
  alias LEFT_BRACKET_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(91);
  alias BACK_SLASH_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(92);
  alias RIGHT_BRACKET_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(93);
  alias HAT_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(94);
  alias UNDERSCORE_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(95);
  alias LEFT_TICK_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(96);
  alias a_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(97);
  alias b_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(98);
  alias c_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(99);
  alias d_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(100);
  alias e_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(101);
  alias f_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(102);
  alias g_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(103);
  alias h_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(104);
  alias i_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(105);
  alias j_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(106);
  alias k_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(107);
  alias l_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(108);
  alias m_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(109);
  alias n_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(110);
  alias o_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(111);
  alias p_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(112);
  alias q_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(113);
  alias r_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(114);
  alias s_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(115);
  alias t_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(116);
  alias u_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(117);
  alias v_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(118);
  alias w_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(119);
  alias x_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(120);
  alias y_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(121);
  alias z_low_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(122);
  alias CURLY_LEFT_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(123);
  alias PIPE_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(124);
  alias CURLY_RIGHT_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(125);
  alias SWUNG_DASH_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(126);
  alias DEL_char: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(127);

end CHARS;