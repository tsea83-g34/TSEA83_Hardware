library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity project is 
    port (clk: std_logic;
          rst: std_logic
    );
end project;

architecture Behavioral of project is 




begin
    process (clk)
    begin
        if rising_edge(clk) then 
            
        end if;




end Behavioral;