library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package PIPECPU_STD is
  
  type byte_mode is (WORD, HALF, BYTE);
  constant PROGRAM_MEMORY_SIZE: INTEGER := 4096;
  constant PROGRAM_MEMORY_ADDRESS_BITS: INTEGER := 12;
  constant PROGRAM_MEMORY_BIT_SIZE: INTEGER := 32;
  constant DATA_MEM_BIT_SIZE: INTEGER := 8;

end PIPECPU_STD;
