library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package CHARS is
  
  constant NUMBER_OF_CHARS : INTEGER := 128;
  constant CHAR_SIZE       : INTEGER := 16;
  
  type char_array is array (0 to NUMBER_OF_CHARS - 1) of UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0);
  
  -- ======== Chars ========
  
  constant CHARS : char_array := (

-- NULL_CHAR
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SOH
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- STX
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ETX
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EOT
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ENQ
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ACK
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- BEL
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- BS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- HT
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- LT
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- VT
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- FF
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- CR
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SO
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SI
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DLE
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DC1
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DC2
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DC3
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DC4
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- NAK
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SYN
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ETB
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- CAN
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EM
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SUB
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ESC
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- FS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- GS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- RS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- US
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SPACE
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EXCLAMATION_MARK
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DOUBLE_QUOTE
"0000000000000000" &
"0000011100111000" &
"0000011100111000" &
"0000011100111000" &
"0000011100111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- HASH
"0000000000000000" &
"0000000011000111" &
"0000000011000111" &
"0000000011000110" &
"0000000011000110" &
"0000111111111111" &
"0000000100001110" &
"0000000100001000" &
"0000000100001000" &
"0011111111111111" &
"0000011000111000" &
"0000011000110000" &
"0000111000110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DOLLAR
"0000000000000000" &
"0000000100000000" &
"0000111111110000" &
"0011100100110000" &
"0011100100000000" &
"1111100100000000" &
"0011111100000000" &
"0000111111110000" &
"0000000111111000" &
"0000000100111000" &
"0000000100111000" &
"0011000100111000" &
"0011111111110000" &
"0000000100000000" &
"0000000100000000" &
"0000000000000000",

-- PERCENT
"0000000000000000" &
"0000000000000000" &
"0000111100000000" &
"0011000011000000" &
"0011000011000000" &
"0011000011000000" &
"0000111100001110" &
"0000000111110000" &
"0000111000111110" &
"0000000011000001" &
"0000000011000001" &
"0000000011000001" &
"0000000000111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- AMPERSAND
"0000000000000000" &
"0000000111110000" &
"0000011000000000" &
"0000011000000000" &
"0000011000000000" &
"0000011100000000" &
"0000111100000000" &
"0000100011000111" &
"0011100011000111" &
"0011100000110111" &
"0011100000001110" &
"0000111000001110" &
"0000011111110111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SINGLE_QUOTE
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- LEFT_PARENTHESES
"0000000000000000" &
"0000000011110000" &
"0000000011000000" &
"0000000111000000" &
"0000000111000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000000111000000" &
"0000000111000000" &
"0000000011000000" &
"0000000011110000" &
"0000000000000000",

-- RIGHT_PARENTHESES
"0000000000000000" &
"0000011100000000" &
"0000000100000000" &
"0000000111000000" &
"0000000111000000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000111000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000000000000000",

-- STAR
"0000000000000000" &
"0000000100000000" &
"0011000100001000" &
"0000100100110000" &
"0000011111000000" &
"0000111111110000" &
"0011000100001000" &
"0000000100000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- PLUS
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111111111110" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- COMMA
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000000000000000",

-- DASH
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- PERIOD
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SLASH
"0000000000000000" &
"0000000000001000" &
"0000000000111000" &
"0000000000110000" &
"0000000011110000" &
"0000000011000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000011000000000" &
"0000111000000000" &
"0000100000000000" &
"0011100000000000" &
"0011100000000000" &
"0000000000000000" &
"0000000000000000",

-- ZERO
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0000100000001000" &
"0011100000001110" &
"0011100000001110" &
"0011100111001110" &
"0011100111001110" &
"0011100000001110" &
"0011100000001110" &
"0000100000001000" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- ONE
"0000000000000000" &
"0000111111000000" &
"0000111111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- TWO
"0000000000000000" &
"0011111111000000" &
"0011000011110000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000011110000" &
"0000000011110000" &
"0000000111000000" &
"0000011100000000" &
"0000111000000000" &
"0011100000000000" &
"0011111111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- THREE
"0000000000000000" &
"0000111111110000" &
"0000000000111110" &
"0000000000001110" &
"0000000000001110" &
"0000000000111000" &
"0000000111000000" &
"0000000000111000" &
"0000000000001110" &
"0000000000001110" &
"0000000000001110" &
"0011000000111000" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- FOUR
"0000000000000000" &
"0000000011111000" &
"0000000011111000" &
"0000000100111000" &
"0000000100111000" &
"0000011000111000" &
"0000111000111000" &
"0000100000111000" &
"0011100000111000" &
"0011111111111111" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- Five
"0000000000000000" &
"0000111111111000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111110000" &
"0000000000111000" &
"0000000000001110" &
"0000000000001110" &
"0000000000001110" &
"0000000000001110" &
"0011000000111000" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SIX
"0000000000000000" &
"0000011111111000" &
"0000111000000000" &
"0000111000000000" &
"0011100000000000" &
"0011100111110000" &
"0011111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SEVEN
"0000000000000000" &
"0011111111111000" &
"0000000000111000" &
"0000000000110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011000000" &
"0000000111000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EIGHT
"0000000000000000" &
"0000011111110000" &
"0011111000111110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- NINE
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111110" &
"0000011111001110" &
"0000000000001110" &
"0000000000111000" &
"0000000000111000" &
"0000111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- COLON
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- SEMICOLON
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000100000000" &
"0000011100000000" &
"0000000000000000",

-- LESS_THAN
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000111" &
"0000000000111110" &
"0000011111110000" &
"0011111000000000" &
"0011111000000000" &
"0000011111110000" &
"0000000000111111" &
"0000000000000110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- EQUAL
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011111111111110" &
"0000000000000000" &
"0000000000000000" &
"0011111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- GREATER_THAN
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011000000000000" &
"0011111100000000" &
"0000000111110000" &
"0000000000001111" &
"0000000000111111" &
"0000000111110000" &
"0011111100000000" &
"0011000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- QUESTION_MARK
"0000000000000000" &
"0000111111110000" &
"0000100000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000011111000" &
"0000000111110000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- AT
"0000000000000000" &
"0000000000000000" &
"0000000111111000" &
"0000011000000110" &
"0000100000000001" &
"0011100011111111" &
"0011000111000111" &
"0011000100000001" &
"0011000100000001" &
"0011000111000111" &
"0011000011111111" &
"0000100000000000" &
"0000100000000000" &
"0000011100000000" &
"0000000111111110" &
"0000000000000000",

-- A
"0000000000000000" &
"0000000111000000" &
"0000011111000000" &
"0000011111110000" &
"0000011011110000" &
"0000011000110000" &
"0000111000110000" &
"0000111000111000" &
"0000100000111000" &
"0011111111111000" &
"0011100000001110" &
"0011000000001110" &
"1111000000000110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- B
"0000000000000000" &
"0011111111110000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011111111000000" &
"0011100000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000111110" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- C
"0000000000000000" &
"0000000111111110" &
"0000111000000110" &
"0000111000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0000111000000000" &
"0000111000000110" &
"0000000111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- D
"0000000000000000" &
"0011111111000000" &
"0011100000111000" &
"0011100000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000111000" &
"0011100000111000" &
"0011111111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- E
"0000000000000000" &
"0000111111111110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111111110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- F
"0000000000000000" &
"0000111111111110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111111110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- G
"0000000000000000" &
"0000000111111000" &
"0000111000001000" &
"0000111000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000" &
"0011100000111110" &
"0011100000001110" &
"0011100000001110" &
"0000100000001110" &
"0000111000001110" &
"0000000111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- H
"0000000000000000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011111111111110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- I
"0000000000000000" &
"0000111111111000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000111111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- J
"0000000000000000" &
"0000011111111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0011000011111000" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- K
"0000000000000000" &
"0011100000001110" &
"0011100000001000" &
"0011100000110000" &
"0011100011110000" &
"0011100111000000" &
"0011111111000000" &
"0011111011000000" &
"0011100011110000" &
"0011100000111000" &
"0011100000111000" &
"0011100000001110" &
"0011100000000111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- L
"0000000000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111111111111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- M
"0000000000000000" &
"0011111000001111" &
"0011111000001111" &
"0011111000001111" &
"0011100100110111" &
"0011100100110111" &
"0011100100110111" &
"0011100011000111" &
"0011100011000111" &
"0011100000000111" &
"0011100000000111" &
"0011100000000111" &
"0011100000000111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- N
"0000000000000000" &
"0011111000001110" &
"0011111000001110" &
"0011111000001110" &
"0011111100001110" &
"0011100100001110" &
"0011100100001110" &
"0011100011001110" &
"0011100011001110" &
"0011100011111110" &
"0011100000111110" &
"0011100000111110" &
"0011100000111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- O
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- P
"0000000000000000" &
"0000111111111000" &
"0000111000001110" &
"0000111000000111" &
"0000111000000111" &
"0000111000000111" &
"0000111000001110" &
"0000111111111000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- Q
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001000" &
"0000111000111000" &
"0000011111110000" &
"0000000000111000" &
"0000000000001000" &
"0000000000000000",

-- R
"0000000000000000" &
"0011111111000000" &
"0011100011110000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100011110000" &
"0011111111000000" &
"0011100011110000" &
"0011100000110000" &
"0011100000001000" &
"0011100000001110" &
"0011100000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- S
"0000000000000000" &
"0000011111111000" &
"0000111000001000" &
"0011100000000000" &
"0011100000000000" &
"0011111000000000" &
"0000111111110000" &
"0000000111111000" &
"0000000000111110" &
"0000000000001110" &
"0000000000001110" &
"0011000000111000" &
"0011111111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- T
"0000000000000000" &
"0011111111111111" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- U
"0000000000000000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- V
"0000000000000000" &
"0011000000001110" &
"0011000000001110" &
"0011100000001000" &
"0011100000001000" &
"0000100000111000" &
"0000100000111000" &
"0000111000110000" &
"0000011000110000" &
"0000011011110000" &
"0000011111110000" &
"0000011111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- W
"0000000000000000" &
"1111000000000111" &
"1111000000000110" &
"1111000000000110" &
"0011000111000110" &
"0011000111000110" &
"0011011111001110" &
"0011011011001110" &
"0011011011111110" &
"0011111000111000" &
"0011111000111000" &
"0000111000111000" &
"0000100000111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- X
"0000000000000000" &
"0011100000001110" &
"0000100000001000" &
"0000111000111000" &
"0000011000110000" &
"0000011111000000" &
"0000000111000000" &
"0000000111000000" &
"0000011111110000" &
"0000111000110000" &
"0000100000111000" &
"0011100000001110" &
"1111000000000110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- Y
"0000000000000000" &
"0011000000000110" &
"0011100000001110" &
"0000100000001000" &
"0000111000111000" &
"0000011111110000" &
"0000011111110000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- Z
"0000000000000000" &
"0011111111111110" &
"0000000000001110" &
"0000000000111000" &
"0000000000110000" &
"0000000011110000" &
"0000000111000000" &
"0000000111000000" &
"0000011100000000" &
"0000011000000000" &
"0000111000000000" &
"0011100000000000" &
"0011111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- LEFT_BRACKET
"0000000000000000" &
"0000000111111000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111111000" &
"0000000000000000",

-- BACK_SLASH
"0000000000000000" &
"0011100000000000" &
"0000100000000000" &
"0000100000000000" &
"0000111000000000" &
"0000011000000000" &
"0000011100000000" &
"0000000100000000" &
"0000000111000000" &
"0000000011000000" &
"0000000011110000" &
"0000000000110000" &
"0000000000111000" &
"0000000000001000" &
"0000000000000000" &
"0000000000000000",

-- RIGHT_BRACKET
"0000000000000000" &
"0000011111110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000000011110000" &
"0000011111110000" &
"0000000000000000",

-- HAT
"0000000000000000" &
"0000000111000000" &
"0000011111110000" &
"0000111000110000" &
"0011100000001000" &
"0011000000000110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- UNDERSCORE
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- LEFT_TICK
"0000011000000000" &
"0000011100000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- a_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111111110000" &
"0000100011111000" &
"0000000000111000" &
"0000000000111000" &
"0000111111111000" &
"0011100000111000" &
"0011100000111000" &
"0011100011111000" &
"0000111100111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- b_low
"0000000000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111011111000" &
"0000111100111000" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111100111000" &
"0000111011111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- c_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000111111110" &
"0000011100000110" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000011100000110" &
"0000000111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- d_low
"0000000000000000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000" &
"0000111100111000" &
"0000111011111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0000111011111000" &
"0000111100111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- e_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011111111111110" &
"0011100000000000" &
"0011100000000000" &
"0000111000000110" &
"0000011111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- f_low
"0000000000000000" &
"0000000011111110" &
"0000000111000000" &
"0000000111000000" &
"0000111111111110" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- g_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111100111000" &
"0000111011111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0000111011111000" &
"0000111100111000" &
"0000000000111000" &
"0000100011110000" &
"0000111111110000",

-- h_low
"0000000000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111011111000" &
"0000111100001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- i_low
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000111111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- j_low
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000000000" &
"0000111111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111100000000",

-- k_low
"0000000000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000000000" &
"0000111000001110" &
"0000111000111000" &
"0000111011110000" &
"0000111111000000" &
"0000111111110000" &
"0000111000111000" &
"0000111000001000" &
"0000111000001110" &
"0000111000000111" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- l_low
"0000000000000000" &
"0000111111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000011111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- m_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011111100111000" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0011100111001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- n_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111011111000" &
"0000111100001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- o_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011111110000" &
"0000111000111000" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0011100000001110" &
"0000111000111000" &
"0000011111110000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- p_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011100111110000" &
"0011111011110000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011111011110000" &
"0011100111110000" &
"0011100000000000" &
"0011100000000000" &
"0011100000000000",

-- q_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111100111000" &
"0000111011111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0011100000111000" &
"0000111011111000" &
"0000111100111000" &
"0000000000111000" &
"0000000000111000" &
"0000000000111000",

-- r_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011100111110" &
"0000011111000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- s_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000011111111000" &
"0000111000000000" &
"0000111000000000" &
"0000111100000000" &
"0000011111111000" &
"0000000000111110" &
"0000000000001110" &
"0000100000001110" &
"0000111111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- t_low
"0000000000000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0011111111111000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000011100000000" &
"0000000111111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- u_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000001110" &
"0000111000111110" &
"0000011111001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- v_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011000000001110" &
"0011100000001000" &
"0000100000111000" &
"0000100000111000" &
"0000111000110000" &
"0000011011110000" &
"0000011011110000" &
"0000011111000000" &
"0000000111000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- w_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"1111000000000111" &
"1111000000000110" &
"0011000000000110" &
"0011000111001110" &
"0011000111001110" &
"0011111011001000" &
"0011111011001000" &
"0000111000111000" &
"0000111000111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- x_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011100000001000" &
"0000111000111000" &
"0000011011110000" &
"0000011111000000" &
"0000000111000000" &
"0000011111000000" &
"0000111000110000" &
"0000100000111000" &
"0011100000001110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- y_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0011000000001000" &
"0011000000111000" &
"0011100000111000" &
"0000100000110000" &
"0000111011110000" &
"0000011011000000" &
"0000011011000000" &
"0000011111000000" &
"0000000100000000" &
"0000011100000000" &
"0000011000000000" &
"0011111000000000",

-- z_low
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111111111110" &
"0000000000001110" &
"0000000000111000" &
"0000000011110000" &
"0000000011000000" &
"0000000111000000" &
"0000011100000000" &
"0000111000000000" &
"0000111111111110" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- CURLY_LEFT
"0000000000000000" &
"0000000011111000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000011111000",

-- PIPE
"0000000000000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000",

-- CURLY_RIGHT
"0000000000000000" &
"0011111100000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000000111000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0000000111000000" &
"0011111100000000",

-- SWUNG_DASH
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000111100000110" &
"0011000011111000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000",

-- DEL
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000" &
"0000000000000000"
);
  
  -- ======== Alias ========
  
  alias NULL_CHAR: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(0);
  alias SOH: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(1);
  alias STX: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(2);
  alias ETX: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(3);
  alias EOT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(4);
  alias ENQ: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(5);
  alias ACK: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(6);
  alias BEL: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(7);
  alias BS: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(8);
  alias HT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(9);
  alias LT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(10);
  alias VT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(11);
  alias FF: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(12);
  alias CR: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(13);
  alias SO: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(14);
  alias SI: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(15);
  alias DLE: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(16);
  alias DC1: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(17);
  alias DC2: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(18);
  alias DC3: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(19);
  alias DC4: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(20);
  alias NAK: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(21);
  alias SYN: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(22);
  alias ETB: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(23);
  alias CAN: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(24);
  alias EM: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(25);
  alias SUB: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(26);
  alias ESC: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(27);
  alias FS: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(28);
  alias GS: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(29);
  alias RS: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(30);
  alias US: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(31);
  alias SPACE: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(32);
  alias EXCLAMATION_MARK: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(33);
  alias DOUBLE_QUOTE: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(34);
  alias HASH: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(35);
  alias DOLLAR: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(36);
  alias PERCENT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(37);
  alias AMPERSAND: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(38);
  alias SINGLE_QUOTE: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(39);
  alias LEFT_PARENTHESES: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(40);
  alias RIGHT_PARENTHESES: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(41);
  alias STAR: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(42);
  alias PLUS: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(43);
  alias COMMA: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(44);
  alias DASH: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(45);
  alias PERIOD: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(46);
  alias SLASH: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(47);
  alias ZERO: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(48);
  alias ONE: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(49);
  alias TWO: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(50);
  alias THREE: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(51);
  alias FOUR: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(52);
  alias Five: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(53);
  alias SIX: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(54);
  alias SEVEN: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(55);
  alias EIGHT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(56);
  alias NINE: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(57);
  alias COLON: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(58);
  alias SEMICOLON: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(59);
  alias LESS_THAN: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(60);
  alias EQUAL: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(61);
  alias GREATER_THAN: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(62);
  alias QUESTION_MARK: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(63);
  alias AT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(64);
  alias A: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(65);
  alias B: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(66);
  alias C: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(67);
  alias D: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(68);
  alias E: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(69);
  alias F: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(70);
  alias G: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(71);
  alias H: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(72);
  alias I: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(73);
  alias J: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(74);
  alias K: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(75);
  alias L: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(76);
  alias M: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(77);
  alias N: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(78);
  alias O: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(79);
  alias P: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(80);
  alias Q: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(81);
  alias R: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(82);
  alias S: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(83);
  alias T: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(84);
  alias U: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(85);
  alias V: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(86);
  alias W: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(87);
  alias X: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(88);
  alias Y: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(89);
  alias Z: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(90);
  alias LEFT_BRACKET: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(91);
  alias BACK_SLASH: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(92);
  alias RIGHT_BRACKET: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(93);
  alias HAT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(94);
  alias UNDERSCORE: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(95);
  alias LEFT_TICK: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(96);
  alias a_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(97);
  alias b_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(98);
  alias c_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(99);
  alias d_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(100);
  alias e_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(101);
  alias f_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(102);
  alias g_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(103);
  alias h_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(104);
  alias i_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(105);
  alias j_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(106);
  alias k_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(107);
  alias l_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(108);
  alias m_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(109);
  alias n_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(110);
  alias o_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(111);
  alias p_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(112);
  alias q_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(113);
  alias r_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(114);
  alias s_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(115);
  alias t_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(116);
  alias u_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(117);
  alias v_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(118);
  alias w_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(119);
  alias x_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(120);
  alias y_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(121);
  alias z_low: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(122);
  alias CURLY_LEFT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(123);
  alias PIPE: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(124);
  alias CURLY_RIGHT: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(125);
  alias SWUNG_DASH: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(126);
  alias DEL: UNSIGNED (CHAR_SIZE * CHAR_SIZE - 1 downto 0) is CHARS(127);

end CHARS;